//----------------------------------------------------------------------
// This File: CYCLE.sv
//----------------------------------------------------------------------
`include "timescale.v"

`ifndef CYCLE_50
  `define CYCLE_50 	20
`endif


`ifndef CYCLE_200
  `define CYCLE_200 5
`endif

`ifndef CYCLE_400
  `define CYCLE_400 2.5
`endif
